*���&O���PH	]�82�xu�z��×���?9����!+�(�gr'-�2���?9H�EExݘ2s�z4p�� (�=8�O��Z��Ue��ħI��`�G/1�{���C0�T�P[���Ws�߮�,c�<A�IM�
uN����"Mϴ-ƛ�dPxD�,!��?/�5PZ��r�L�����pyт�O�1�6���@42�>N�I�N��;��>z���|Dd>;�N��q �XECÀ����u?�ʒ��\�B; � ��LX3<qu�<���R�l�}V@�L(����yUl|\>� o<|}>�΂P6	@aʁ@���m1��L,��М�F4k�*��